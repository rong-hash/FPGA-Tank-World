module coin_silver_rom (
	input logic clock,
	input logic [12:0] address,
	output logic [1:0] q
);

logic [1:0] memory [0:8191] /* synthesis ram_init_file = "./coin_silver/coin_silver.mif" */;

always_ff @ (posedge clock) begin
	q <= memory[address];
end

endmodule
